module IntToSeg(

);
