module Starter(
          input Clk100M,
          input ,
          output start,
);

endmodule