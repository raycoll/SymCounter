///////////////////////////////////
// Outputs a signal to 
///////////////////////////////////
module CurPeriod(
          input Clk100M,
          input prelimSig,
          input gameSig,
          input answerSig,
          input postSig,
          output reg pre,
          output reg game,
          output reg answer,
          output reg post
);


endmodule