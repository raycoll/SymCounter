module SymGen(
                input 
);