module PrelimPeriod(
          input Clk1Hz,
          input prelimSig,
          output gameSig,
          output reg [7:0] prelimSeg0,
          output reg [7:0] prelimSeg1,
          output reg [7:0] prelimSeg2,
          output reg [7:0] prelimSeg3
);

