module DispCntrl(
                
);